// YARP UVM Package - Top-level package that includes all verification components
package yarp_uvm_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  import yarp_pkg::*;
  import yarp_seq_pkg::*;
  import yarp_agent_pkg::*;
  import yarp_env_pkg::*;
  import yarp_test_pkg::*;
  
endpackage
